LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE ULA_PACKAGE IS

	COMPONENT DECODIFICADOR_3x8 IS
		PORT(SEL: BIT_VECTOR (2 DOWNTO 0);
			 S : OUT BIT_VECTOR(7 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT DECODIFICADOR_8X1 IS
		PORT(SEL: BIT_VECTOR (2 DOWNTO 0);
			 S : OUT BIT_VECTOR(7 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT PORTAS_LOGICAS IS
		PORT(A,B: IN BIT;
			 E_PL: IN BIT_VECTOR;
			 S: OUT BIT_VECTOR(5 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT SOMADOR IS
		PORT (A_B_Cin: IN BIT_VECTOR (2 DOWNTO 0);    
		      S_Cout: OUT BIT_vector (1 DOWNTO 0));
	END COMPONENT;

	COMPONENT SUBTRATOR IS
		PORT(EN_SUB: IN BIT_VECTOR (2 DOWNTO 0);
		     S_Cout: OUT BIT_VECTOR (1 DOWNTO 0));
	END COMPONENT;

END ULA_PACKAGE;