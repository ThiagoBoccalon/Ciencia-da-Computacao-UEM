LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE DECODIFICADOR_PACKAGE IS
	
	COMPONENT NOT_1 IS
		PORT(A: IN BIT;
		 S: OUT BIT);
	END COMPONENT;

	COMPONENT AND_2 IS
		PORT(A,B: IN BIT;
		 S: OUT BIT);
	END COMPONENT;

END DECODIFICADOR_PACKAGE;

ENTITY DECODIFICADOR IS
	PORT(EN_DC: IN BIT_VECTOR (2 DOWNTO 0);
		 S_UL0, S_UL1: OUT BIT;
		 S_PC0, S_PC1, S_PC2, S_PC3, S_PC4, S_PC5: OUT BIT); -- S_UL S�O AS SAIDAS PARA AS UNIDADES L�GICAS DA ULA
																				 -- J� AS SAIDA S_PC S�O SAIDAS PARA AS PORTAS DE CONTROLE DA ULA	
END DECODIFICADOR;

ARCHITECTURE TEST_DECODIFICADOR OF DECODIFICADOR IS
BEGIN
		PROCESS(EN_DC)
		BEGIN
				CASE EN_DC IS
					WHEN "000" => S_PC5 <= '1';
					WHEN "001" => S_PC4 <= '1';
					WHEN "010" => S_PC3 <= '1';
					WHEN "011" => S_PC2 <= '1';
					WHEN "100" => S_PC1 <= '1';
					WHEN "101" => S_PC0 <= '1';
					WHEN "110" => S_UL0 <= '1';
					WHEN "111" => S_UL1 <= '1';
				END CASE;
		END PROCESS;
END TEST_DECODIFICADOR;