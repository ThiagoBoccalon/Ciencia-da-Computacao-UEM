LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE MUX_2X1_PACKAGE IS
	
	COMPONENT NOT_1 IS
		PORT(A: IN BIT;
			 Z: OUT BIT);
	END COMPONENT;
	
	COMPONENT AND_2 IS 
		PORT(A,B: IN BIT;
			 Z: OUT BIT);
	END COMPONENT;
	
	COMPONENT OR_2 IS
		PORT(A,B: IN BIT;
		     Z: OUT BIT);
	END COMPONENT;
	
END MUX_2X1_PACKAGE;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

	-- PACOTE
	
	USE WORK_2.MUX_2X1_PACKAGE.ALL;
	
	-- DECLARA ENTIDADE PARA O PACOTE DE MUX 2X1

ENTITY MUX_2X1 IS
	PORT(S0,S1,CH: IN BIT;
		 F: OUT BIT);
END MUX_2X1;


ARCHITECTURE ESTRUTURAL OF MUX_2X1 IS
	
	SIGNAL T0, T1, T2: BIT;
	
BEGIN 
	P1: NOT_1 PORT MAP (CH,T0);
	P2: AND_2 PORT MAP (S0,T0,T1);
	P3: AND_2 PORT MAP (CH,S1,T2);
	P4: OR_2 PORT MAP (T1,T2,F);
END ESTRUTURAL;
	
	
	



	