LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY AND_3 IS
	PORT(A,B,C: IN BIT;
		 S: OUT BIT);
END AND_3;

ARCHITECTURE TEST_2 OF AND_3 IS
BEGIN
	S <= A AND B AND 3;
END TEST_2;