library ieee;
use ieee.std_logic_1164.all;

Entity Exercicio_1_Case_When is
	Port ( Re, Vre, Asg, Sct: 
			) -- 