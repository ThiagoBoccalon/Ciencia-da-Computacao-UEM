LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REL_SEG_MIN IS
	PORT(CLK,RST: IN BIT;
		  )
END REL_SEG_MIN;

ARCHITECTURE ESTRUTURAL OF IS

SIGNAL LEVA: 

COMPONENT CONT_SEG IS
	PORT(CLK, RST: IN BIT;
		 RCO: OUT BIT;
		 UNID, DEZ: OUT INTEGER RANGE 0 TO 15);
END COMPONENT;

BEGIN
	P_MIN: 