LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FFD_C is
	PORT(CLR, CLK, D: IN STD_LOGIC;
		 Q, QBAR: BUFFER STD_LOGIC);
END FFD_C;

ARCHITECTURE COMPORTAMENTAL OF FFD_C IS
BEGIN
	PROCESS(CLR,CLK,D)
	VARIABLE QV, QBARV: STD_LOGIC;
	BEGIN
	IF (CLR ='0') THEN
		QV:= '0';
		QBARV:= NOT QV;
	ELSIF (FALLING_EDGE(CLK)) THEN
		QV:= D;
		QBARV:= NOT D;
	END IF;
	Q <= QV;
	QBAR <= NOT Q;
	END PROCESS;
END COMPORTAMENTAL;