LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY OR_8 IS
	PORT(A,B,C,D,E,F,G,H: IN BIT;
		 S: OUT BIT);
END OR_8;

ARCHITECTURE TEST_OR OF OR_8 IS
BEGIN
		S <= A OR B OR C OR D OR E OR F OR G OR H;
END TEST_OR;