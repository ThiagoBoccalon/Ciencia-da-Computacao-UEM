LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY OR_2 IS
	PORT(A,B: IN BIT;
		 Z: OUT BIT);
END OR_2;

ARCHITECTURE TEST3 OF OR_2 IS 
	BEGIN
		Z <= A OR B;
	END TEST3;