CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 4 110 10
176 75 1278 973
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 171 457 268
9437202 0
0
6 Title:
5 Name:
0
0
0
7
7 Ground~
168 36 395 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5130 0 0
2
39614.8 1
0
7 Pulser~
4 310 405 0 10 12
0 17 18 7 19 0 0 10 10 8
8
0
0 0 4656 512
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
391 0 0
2
39614.8 0
0
2 +V
167 29 47 0 1 3
0 6
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3124 0 0
2
39614.8 0
0
9 CA 7-Seg~
184 173 124 0 18 19
10 14 13 12 11 10 9 8 20 6
2 0 0 2 2 0 0 2 1
0
0 0 21088 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
3421 0 0
2
39614.8 0
0
6 74LS47
187 181 223 0 14 29
0 16 5 4 15 6 21 8 9 10
11 12 13 14 6
0
0 0 4848 90
7 74LS247
-24 -60 25 -52
2 U3
60 0 74 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 0 0 0 0
1 U
8157 0 0
2
39614.8 0
0
6 74LS90
107 173 338 0 10 21
0 2 2 3 3 7 15 16 5 4
15
0
0 0 4848 90
6 74LS90
-21 -51 21 -43
2 U2
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 0 0 0 0
1 U
5572 0 0
2
39614.8 0
0
9 2-In AND~
219 66 283 0 3 22
0 4 5 3
0
0 0 624 512
5 74F08
-18 -24 17 -16
3 U1A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
8901 0 0
2
39614.8 0
0
24
0 4 3 0 0 4096 0 0 6 2 0 3
163 373
173 373
173 364
3 3 3 0 0 8320 0 7 6 0 0 4
41 283
41 373
164 373
164 364
2 0 2 0 0 4096 0 6 0 0 5 2
155 364
155 389
1 0 2 0 0 0 0 6 0 0 5 2
146 364
146 389
1 0 2 0 0 4224 0 1 0 0 0 2
36 389
173 389
1 0 4 0 0 8320 0 7 0 0 21 3
86 274
86 273
165 273
0 2 5 0 0 8320 0 0 7 20 0 3
155 291
155 292
86 292
5 0 6 0 0 12288 0 5 0 0 24 4
218 260
218 264
272 264
272 56
14 0 6 0 0 0 0 5 0 0 24 4
227 196
227 61
228 61
228 56
5 3 7 0 0 8320 0 6 2 0 0 3
191 370
191 396
286 396
7 7 8 0 0 8320 0 5 4 0 0 4
146 190
146 183
188 183
188 160
8 6 9 0 0 8320 0 5 4 0 0 4
155 190
155 183
182 183
182 160
9 5 10 0 0 12416 0 5 4 0 0 4
164 190
164 183
176 183
176 160
10 4 11 0 0 12416 0 5 4 0 0 4
173 190
173 183
170 183
170 160
11 3 12 0 0 8320 0 5 4 0 0 4
182 190
182 178
164 178
164 160
12 2 13 0 0 8320 0 5 4 0 0 4
191 190
191 173
158 173
158 160
13 1 14 0 0 8320 0 5 4 0 0 4
200 190
200 168
152 168
152 160
6 10 15 0 0 12416 0 6 6 0 0 6
200 370
200 374
215 374
215 292
200 292
200 300
1 7 16 0 0 4224 0 5 6 0 0 2
146 260
146 300
2 8 5 0 0 128 0 5 6 0 0 4
155 260
155 292
164 292
164 300
9 3 4 0 0 128 0 6 5 0 0 4
182 300
182 273
164 273
164 260
10 4 15 0 0 0 0 6 5 0 0 4
200 300
200 268
173 268
173 260
9 0 6 0 0 0 0 4 0 0 24 2
173 88
173 56
1 0 6 0 0 4224 0 3 0 0 0 3
29 56
878 56
878 66
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
