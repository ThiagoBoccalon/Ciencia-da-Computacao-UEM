-- SOMADOR COMPLETO DE 1 BIT
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SOMADOR IS
	PORT (A_B_Cin: IN BIT_VECTOR (2 downTO 0);   -- A = (2), B(1), Cin(0)
		  S_Cout: OUT BIT_vector (1 downto 0)); -- DA UMA VERIFICADA AQUI MAS ACHO QUE � S� 1 BIT QUE SAI
END SOMADOR;

-- O SOMADOR DEVE SER FEITO USANDO WHITE SELECT WHEN

ARCHITECTURE TEST_SOMADOR OF SOMADOR IS
	BEGIN
		WITH A_B_Cin SELECT
			S_Cout <= "00" WHEN "000",
				      "10" WHEN "001",
				      "10" WHEN "010",
				      "01" WHEN "011",
				      "10" WHEN "100",
				      "01" WHEN "101",
				      "01" WHEN "110",
				      "11" WHEN "111";
	END TEST_SOMADOR;