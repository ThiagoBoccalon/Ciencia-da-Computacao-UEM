LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY EXERCICIO_9_SELECT_WHEN IS
	PORT( CH: IN BIT_VECTOR (2 DOWNTO 0);
	      S1: OUT BIT_VECTOR (3 DOWNTO 0));
END EXERCICIO_9_SELECT_WHEN;

ARCHITECTURE TEST OF EXERCICIO_9_SELECT_WHEN IS
BEGIN
	WITH CH SELECT
		S1 <= "0000" WHEN "000" | "010" | "100" | "110",
			  "1000" WHEN "001",
			  "0010" WHEN "011",
			  "0100" WHEN "101",
			  "0001" WHEN "111";
END TEST; 	 