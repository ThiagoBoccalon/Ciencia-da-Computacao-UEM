LIBRARY IEEE;
IEEE.STD_LOGIC_1164.ALL;

ENTITY DECODIFICADOR_8x1 IS 
	PORT(SEL: BIT_VECTOR (2 DOWNTO 0);
		 E_SOM, E_SUB, E3, E4, E5, E6, E7, E8: IN BIT;	
		 SAIDA_ULA: OUT BIT);
ENTITY DECODIFICADOR_8x1;

ARCHITECTURE TEST_DECO_8x1 OF DECODIFICADOR_8x1 IS
	BEGIN
		PROCESS(SEL)
			BEGIN
				CASE SEL IS
					WHEN "000" => SAIDA_ULA <= "E_SOM"; 
					WHEN "001" => SAIDA_ULA <= "E_SUB";
					WHEN "010" => SAIDA_ULA <= "E3";
					WHEN "011" => SAIDA_ULA <= "E4";
					WHEN "100" => SAIDA_ULA <= "E5";
					WHEN "101" => SAIDA_ULA <= "E6";
					WHEN "110" => SAIDA_ULA <= "E7"; 
					WHEN "111" => SAIDA_ULA <= "E8"; 
				END CASE;