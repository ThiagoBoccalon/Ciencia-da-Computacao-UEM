CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 77 1438 849
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 173 457 270
9437202 0
0
6 Title:
5 Name:
0
0
0
27
9 2-In AND~
219 179 362 0 3 22
0 4 3 5
0
0 0 624 782
6 74LS08
-21 -24 21 -16
4 U14B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
5130 0 0
2
39570.9 0
0
9 2-In AND~
219 169 506 0 3 22
0 9 8 7
0
0 0 624 512
6 74LS08
-21 -24 21 -16
4 U14A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
391 0 0
2
5.89388e-315 0
0
9 2-In AND~
219 290 511 0 3 22
0 11 10 6
0
0 0 624 512
6 74LS08
-21 -24 21 -16
4 U13D
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3124 0 0
2
5.89388e-315 0
0
9 2-In AND~
219 490 534 0 3 22
0 13 14 12
0
0 0 624 512
6 74LS08
-21 -24 21 -16
4 U13C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3421 0 0
2
5.89388e-315 0
0
9 2-In AND~
219 650 559 0 3 22
0 16 17 15
0
0 0 624 692
6 74LS08
-21 -24 21 -16
4 U13B
-17 -25 11 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
8157 0 0
2
5.89388e-315 0
0
9 2-In AND~
219 756 498 0 3 22
0 19 20 18
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U13A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5572 0 0
2
39570.9 0
0
7 Pulser~
4 937 489 0 10 12
0 77 78 67 79 0 0 1 1 1
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8901 0 0
2
5.89388e-315 0
0
7 Ground~
168 51 454 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
5.89388e-315 5.26354e-315
0
6 74LS47
187 837 232 0 14 29
0 20 68 69 19 80 81 60 61 62
63 64 65 66 24
0
0 0 4848 90
7 74LS247
-24 -60 25 -52
3 U11
59 0 80 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4747 0 0
2
5.89388e-315 5.30499e-315
0
9 CA 7-Seg~
184 825 110 0 18 19
10 66 65 64 63 62 61 60 82 24
2 0 0 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP5
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
972 0 0
2
5.89388e-315 5.32571e-315
0
6 74LS47
187 104 225 0 14 29
0 75 76 4 21 83 84 53 54 55
56 57 58 59 24
0
0 0 4848 90
7 74LS247
-24 -60 25 -52
3 U12
59 0 80 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3472 0 0
2
5.89388e-315 5.34643e-315
0
9 CA 7-Seg~
184 92 103 0 18 19
10 59 58 57 56 55 54 53 85 24
0 0 0 0 0 0 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP6
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9998 0 0
2
5.89388e-315 5.3568e-315
0
9 CA 7-Seg~
184 239 103 0 18 19
10 52 51 50 49 48 47 46 86 24
2 0 0 2 2 2 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3536 0 0
2
5.89388e-315 5.36716e-315
0
6 74LS47
187 251 225 0 14 29
0 9 3 74 8 87 88 46 47 48
49 50 51 52 24
0
0 0 4848 90
7 74LS247
-24 -60 25 -52
2 U7
62 0 76 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
4597 0 0
2
5.89388e-315 5.37752e-315
0
9 CA 7-Seg~
184 391 104 0 18 19
10 45 44 43 42 41 40 39 89 24
0 0 0 0 0 0 2 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3835 0 0
2
5.89388e-315 5.38788e-315
0
6 74LS47
187 403 226 0 14 29
0 73 11 10 22 90 91 39 40 41
42 43 44 45 24
0
0 0 4848 90
7 74LS247
-24 -60 25 -52
2 U8
62 0 76 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3670 0 0
2
5.89388e-315 5.39306e-315
0
9 CA 7-Seg~
184 537 108 0 18 19
10 38 37 36 35 34 33 32 92 24
0 2 0 0 2 0 0 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
5616 0 0
2
5.89388e-315 5.39824e-315
0
6 74LS47
187 549 230 0 14 29
0 14 71 72 13 93 94 32 33 34
35 36 37 38 24
0
0 0 4848 90
7 74LS247
-24 -60 25 -52
2 U9
62 0 76 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
9323 0 0
2
5.89388e-315 5.40342e-315
0
9 CA 7-Seg~
184 678 110 0 18 19
10 31 30 29 28 27 26 25 95 24
0 0 2 0 0 2 0 2 1
0
0 0 21104 0
5 REDCA
16 -41 51 -33
5 DISP4
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
317 0 0
2
5.89388e-315 5.4086e-315
0
6 74LS47
187 690 232 0 14 29
0 70 17 16 23 96 97 25 26 27
28 29 30 31 24
0
0 0 4848 90
7 74LS247
-24 -60 25 -52
3 U10
59 0 80 8
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3108 0 0
2
5.89388e-315 5.41378e-315
0
2 +V
167 13 28 0 1 3
0 24
0
0 0 54256 0
2 5v
-8 -22 6 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4299 0 0
2
5.89388e-315 5.41896e-315
0
6 74LS90
107 108 387 0 10 21
0 2 2 5 5 7 21 75 76 4
21
0
0 0 4848 90
6 74LS90
-21 -51 21 -43
2 U6
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
9672 0 0
2
5.89388e-315 5.42414e-315
0
6 74LS90
107 246 389 0 10 21
0 2 2 5 5 6 8 9 3 74
8
0
0 0 4848 90
6 74LS90
-21 -51 21 -43
2 U5
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
7876 0 0
2
5.89388e-315 5.42933e-315
0
6 74LS90
107 396 393 0 10 21
0 2 2 6 6 12 22 73 11 10
22
0
0 0 4848 90
6 74LS90
-21 -51 21 -43
2 U4
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
6369 0 0
2
5.89388e-315 5.43192e-315
0
6 74LS90
107 544 392 0 10 21
0 2 2 2 2 15 13 14 71 72
13
0
0 0 4848 90
6 74LS90
-21 -51 21 -43
2 U3
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
9172 0 0
2
5.89388e-315 5.43451e-315
0
6 74LS90
107 689 396 0 10 21
0 2 2 15 15 18 23 70 17 16
23
0
0 0 4848 90
6 74LS90
-21 -51 21 -43
2 U2
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
7100 0 0
2
5.89388e-315 5.4371e-315
0
6 74LS90
107 845 395 0 10 21
0 2 2 2 2 67 19 20 68 69
19
0
0 0 4848 90
6 74LS90
-21 -51 21 -43
2 U1
41 -11 55 -3
0
15 DVCC=5;DGND=10;
93 %D [%5bi %10bi %1i %2i %3i %4i %5i %6i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o] %M
0
12 type:digital
5 DIP14
21

0 6 7 2 3 14 1 11 8 9
12 6 7 2 3 14 1 11 8 9
12 0
65 0 0 0 1 0 0 0
1 U
3820 0 0
2
5.89388e-315 5.43969e-315
0
127
2 0 3 0 0 4096 0 1 0 0 114 3
186 340
186 287
237 287
1 0 4 0 0 4096 0 1 0 0 119 3
168 340
168 275
117 275
3 0 2 0 0 4096 0 25 0 0 96 2
535 418
535 440
4 0 2 0 0 0 0 25 0 0 96 2
544 418
544 440
4 0 5 0 0 4096 0 23 0 0 6 4
246 415
246 430
236 430
236 427
0 3 5 0 0 4096 0 0 23 8 0 3
180 427
237 427
237 415
0 3 5 0 0 0 0 0 22 8 0 3
108 427
99 427
99 413
3 4 5 0 0 16512 0 1 22 0 0 6
177 385
177 427
180 427
180 427
108 427
108 413
0 4 6 0 0 8192 0 0 24 10 0 3
387 453
396 453
396 419
0 3 6 0 0 4224 0 0 24 14 0 3
264 467
387 467
387 419
3 5 7 0 0 8320 0 2 22 0 0 3
144 506
126 506
126 419
0 2 8 0 0 8320 0 0 2 116 0 4
273 346
198 346
198 515
189 515
0 1 9 0 0 8320 0 0 2 113 0 4
219 347
198 347
198 497
189 497
3 5 6 0 0 0 0 3 23 0 0 3
265 511
264 511
264 421
0 2 10 0 0 8320 0 0 3 111 0 4
405 345
322 345
322 520
310 520
0 1 11 0 0 8320 0 0 3 110 0 4
387 346
325 346
325 502
310 502
3 5 12 0 0 8320 0 4 24 0 0 3
465 534
414 534
414 425
0 1 13 0 0 8320 0 0 4 108 0 6
571 348
473 348
473 459
544 459
544 525
510 525
0 2 14 0 0 8320 0 0 4 105 0 6
514 350
483 350
483 485
539 485
539 543
510 543
0 5 15 0 0 8192 0 0 25 22 0 4
689 489
689 482
562 482
562 424
3 3 15 0 0 0 0 5 26 0 0 5
671 559
682 559
682 436
680 436
680 422
3 4 15 0 0 8320 0 5 26 0 0 3
671 559
689 559
689 422
0 1 16 0 0 8320 0 0 5 103 0 4
698 351
620 351
620 568
626 568
0 2 17 0 0 12416 0 0 5 102 0 5
680 349
680 354
625 354
625 550
626 550
3 5 18 0 0 8320 0 6 26 0 0 3
729 498
707 498
707 428
0 1 19 0 0 8320 0 0 6 100 0 4
872 348
789 348
789 507
774 507
0 2 20 0 0 8320 0 0 6 97 0 4
802 343
784 343
784 489
774 489
6 0 19 0 0 0 0 27 0 0 100 5
872 427
872 431
887 431
887 315
872 315
2 0 2 0 0 0 0 26 0 0 96 2
671 422
671 440
1 0 2 0 0 0 0 26 0 0 96 2
662 422
662 440
6 0 21 0 0 12416 0 22 0 0 120 5
135 419
135 423
150 423
150 326
135 326
6 0 8 0 0 0 0 23 0 0 116 5
273 421
273 425
288 425
288 327
273 327
6 0 22 0 0 12416 0 24 0 0 112 5
423 425
423 429
438 429
438 322
423 322
6 0 13 0 0 0 0 25 0 0 108 5
571 424
571 428
586 428
586 327
571 327
6 0 23 0 0 12416 0 26 0 0 104 5
716 428
716 431
731 431
731 327
716 327
0 9 24 0 0 4096 0 0 19 127 0 2
678 37
678 74
7 7 25 0 0 8320 0 20 19 0 0 4
655 199
655 179
693 179
693 146
8 6 26 0 0 12416 0 20 19 0 0 4
664 199
664 174
687 174
687 146
9 5 27 0 0 4224 0 20 19 0 0 4
673 199
673 169
681 169
681 146
10 4 28 0 0 4224 0 20 19 0 0 4
682 199
682 164
675 164
675 146
11 3 29 0 0 4224 0 20 19 0 0 4
691 199
691 159
669 159
669 146
2 12 30 0 0 4224 0 19 20 0 0 4
663 146
663 191
700 191
700 199
13 1 31 0 0 8320 0 20 19 0 0 4
709 199
709 154
657 154
657 146
0 9 24 0 0 0 0 0 17 127 0 2
537 37
537 72
7 7 32 0 0 8320 0 18 17 0 0 4
514 197
514 177
552 177
552 144
8 6 33 0 0 12416 0 18 17 0 0 4
523 197
523 172
546 172
546 144
9 5 34 0 0 4224 0 18 17 0 0 4
532 197
532 167
540 167
540 144
10 4 35 0 0 4224 0 18 17 0 0 4
541 197
541 162
534 162
534 144
11 3 36 0 0 4224 0 18 17 0 0 4
550 197
550 157
528 157
528 144
2 12 37 0 0 4224 0 17 18 0 0 4
522 144
522 189
559 189
559 197
13 1 38 0 0 8320 0 18 17 0 0 4
568 197
568 152
516 152
516 144
0 9 24 0 0 0 0 0 15 127 0 2
391 37
391 68
7 7 39 0 0 8320 0 16 15 0 0 4
368 193
368 173
406 173
406 140
8 6 40 0 0 12416 0 16 15 0 0 4
377 193
377 168
400 168
400 140
9 5 41 0 0 4224 0 16 15 0 0 4
386 193
386 163
394 163
394 140
10 4 42 0 0 4224 0 16 15 0 0 4
395 193
395 158
388 158
388 140
11 3 43 0 0 4224 0 16 15 0 0 4
404 193
404 153
382 153
382 140
2 12 44 0 0 4224 0 15 16 0 0 4
376 140
376 185
413 185
413 193
13 1 45 0 0 8320 0 16 15 0 0 4
422 193
422 148
370 148
370 140
0 9 24 0 0 0 0 0 13 127 0 2
239 37
239 67
7 7 46 0 0 8320 0 14 13 0 0 4
216 192
216 172
254 172
254 139
8 6 47 0 0 12416 0 14 13 0 0 4
225 192
225 167
248 167
248 139
9 5 48 0 0 4224 0 14 13 0 0 4
234 192
234 162
242 162
242 139
10 4 49 0 0 4224 0 14 13 0 0 4
243 192
243 157
236 157
236 139
11 3 50 0 0 4224 0 14 13 0 0 4
252 192
252 152
230 152
230 139
2 12 51 0 0 4224 0 13 14 0 0 4
224 139
224 184
261 184
261 192
13 1 52 0 0 8320 0 14 13 0 0 4
270 192
270 147
218 147
218 139
0 9 24 0 0 0 0 0 12 127 0 2
92 37
92 67
7 7 53 0 0 8320 0 11 12 0 0 4
69 192
69 172
107 172
107 139
8 6 54 0 0 12416 0 11 12 0 0 4
78 192
78 167
101 167
101 139
9 5 55 0 0 4224 0 11 12 0 0 4
87 192
87 162
95 162
95 139
10 4 56 0 0 4224 0 11 12 0 0 4
96 192
96 157
89 157
89 139
11 3 57 0 0 4224 0 11 12 0 0 4
105 192
105 152
83 152
83 139
2 12 58 0 0 4224 0 12 11 0 0 4
77 139
77 184
114 184
114 192
13 1 59 0 0 8320 0 11 12 0 0 4
123 192
123 147
71 147
71 139
0 9 24 0 0 0 0 0 10 127 0 2
825 37
825 74
7 7 60 0 0 8320 0 9 10 0 0 4
802 199
802 179
840 179
840 146
8 6 61 0 0 12416 0 9 10 0 0 4
811 199
811 174
834 174
834 146
9 5 62 0 0 4224 0 9 10 0 0 4
820 199
820 169
828 169
828 146
10 4 63 0 0 4224 0 9 10 0 0 4
829 199
829 164
822 164
822 146
11 3 64 0 0 4224 0 9 10 0 0 4
838 199
838 159
816 159
816 146
2 12 65 0 0 4224 0 10 9 0 0 4
810 146
810 191
847 191
847 199
13 1 66 0 0 8320 0 9 10 0 0 4
856 199
856 154
804 154
804 146
5 3 67 0 0 8320 0 27 7 0 0 5
863 427
863 466
975 466
975 480
961 480
3 0 2 0 0 0 0 27 0 0 96 2
836 421
836 440
2 0 2 0 0 0 0 27 0 0 96 2
827 421
827 440
1 0 2 0 0 0 0 27 0 0 96 2
818 421
818 440
2 0 2 0 0 0 0 25 0 0 96 2
526 418
526 440
1 0 2 0 0 0 0 25 0 0 96 2
517 418
517 440
2 0 2 0 0 0 0 24 0 0 96 2
378 419
378 440
1 0 2 0 0 0 0 24 0 0 96 2
369 419
369 440
2 0 2 0 0 4096 0 23 0 0 96 2
228 415
228 440
1 0 2 0 0 0 0 23 0 0 96 2
219 415
219 440
2 0 2 0 0 4096 0 22 0 0 96 2
90 413
90 440
1 0 2 0 0 0 0 22 0 0 96 2
81 413
81 440
1 4 2 0 0 8320 0 8 27 0 0 4
51 448
51 440
845 440
845 421
1 7 20 0 0 0 0 9 27 0 0 4
802 269
802 344
818 344
818 357
2 8 68 0 0 4224 0 9 27 0 0 4
811 269
811 349
836 349
836 357
9 3 69 0 0 4224 0 27 9 0 0 4
854 357
854 282
820 282
820 269
10 4 19 0 0 0 0 27 9 0 0 4
872 357
872 277
829 277
829 269
1 7 70 0 0 4224 0 20 26 0 0 4
655 269
655 349
662 349
662 358
2 8 17 0 0 0 0 20 26 0 0 4
664 269
664 349
680 349
680 358
9 3 16 0 0 0 0 26 20 0 0 4
698 358
698 282
673 282
673 269
10 4 23 0 0 0 0 26 20 0 0 4
716 358
716 277
682 277
682 269
1 7 14 0 0 0 0 18 25 0 0 4
514 267
514 346
517 346
517 354
2 8 71 0 0 4224 0 18 25 0 0 4
523 267
523 346
535 346
535 354
9 3 72 0 0 4224 0 25 18 0 0 4
553 354
553 280
532 280
532 267
10 4 13 0 0 0 0 25 18 0 0 4
571 354
571 275
541 275
541 267
1 7 73 0 0 4224 0 16 24 0 0 4
368 263
368 347
369 347
369 355
8 2 11 0 0 0 0 24 16 0 0 4
387 355
387 271
377 271
377 263
9 3 10 0 0 0 0 24 16 0 0 4
405 355
405 276
386 276
386 263
10 4 22 0 0 0 0 24 16 0 0 4
423 355
423 271
395 271
395 263
7 1 9 0 0 0 0 23 14 0 0 4
219 351
219 270
216 270
216 262
8 2 3 0 0 4224 0 23 14 0 0 4
237 351
237 270
225 270
225 262
9 3 74 0 0 4224 0 23 14 0 0 4
255 351
255 275
234 275
234 262
10 4 8 0 0 0 0 23 14 0 0 4
273 351
273 270
243 270
243 262
7 1 75 0 0 4224 0 22 11 0 0 4
81 349
81 291
69 291
69 262
8 2 76 0 0 4224 0 22 11 0 0 4
99 349
99 280
78 280
78 262
9 3 4 0 0 4224 0 22 11 0 0 4
117 349
117 275
87 275
87 262
10 4 21 0 0 0 0 22 11 0 0 4
135 349
135 270
96 270
96 262
14 0 24 0 0 4096 0 9 0 0 127 2
883 205
883 37
14 0 24 0 0 0 0 20 0 0 127 2
736 205
736 37
14 0 24 0 0 0 0 18 0 0 127 2
595 203
595 37
14 0 24 0 0 0 0 16 0 0 127 2
449 199
449 37
14 0 24 0 0 0 0 14 0 0 127 2
297 198
297 37
14 0 24 0 0 0 0 11 0 0 127 2
150 198
150 37
1 0 24 0 0 4224 0 21 0 0 0 2
13 37
917 37
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 5e-06 2e-08 2e-08
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
