Library ieee;
Use ieee.std_logic_1164.all; -- nesse pacote est�o todos os componentes utilizados
Package blocos_package is
COMPONENT PORTAS_LOGICAS IS
	PORT(A_B_Cin : IN BIT_VECTOR (2 DOWNTO 0);
		Saida_deco : IN BIT_VECTOR (7 DOWNTO 0);
		S: OUT BIT);
END COMPONENT;
COMPONENT SELECAO_SAIDA IS
	PORT( S_SOM,S_SUB,Cout_SOM,Cout_SUB,S_LOGICA : IN BIT;
		  S,Cout : OUT BIT); 
END COMPONENT;
COMPONENT SOMADOR IS
	PORT (A_B_Cin: IN BIT_VECTOR (2 DOWNTO 0);
		  SAIDA_DECO : IN BIT_VECTOR(7 DOWNTO 0);		      
		  S_SOM, Cout_SOM: OUT BIT;
		  S,Cout: BUFFER BIT);
END COMPONENT;

COMPONENT SUBTRATOR IS
	PORT(EN_SUB: IN BIT_VECTOR (2 DOWNTO 0);
		 SAIDA_DECO : IN BIT_VECTOR(7 DOWNTO 0);
		 S_SUB,Cout_SUB : OUT BIT;
		 S,Cout: BUFFER BIT);
END COMPONENT;

COMPONENT DECODIFICADOR_3X8 IS
	PORT(SEL: BIT_VECTOR (2 DOWNTO 0);
		 S : OUT BIT_VECTOR(7 DOWNTO 0));
END COMPONENT;
end blocos_package;