LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY PORTAS_LOGICAS IS
	PORT(A_B_Cin : IN BIT_VECTOR (2 DOWNTO 0);
		Saida_deco : IN BIT_VECTOR (7 DOWNTO 0);
		S_Cout, S_Cout2 : IN BIT_VECTOR (1 DOWNTO 0);
		S, Cout: OUT BIT);
END PORTAS_LOGICAS;
ARCHITECTURE COMPORTAMENTAL OF PORTAS_LOGICAS IS
BEGIN
		PROCESS(A_B_Cin, saida_deco, S_Cout, S_Cout2)
		BEGIN	
			Cout <= '0';
			IF (saida_deco(0)= '1') THEN
				S <= A_B_Cin(2) AND A_B_Cin(1); -- s0 estar� recebendo A e B
			ELSIF (saida_deco(1)= '1') THEN
				S <= A_B_Cin(2) NAND A_B_Cin(1);
			ELSIF (saida_deco(2)= '1') THEN
				S <= A_B_Cin(2) OR A_B_Cin(1);
			ELSIF (saida_deco(3)= '1') THEN
				S <= A_B_Cin(2) NOR A_B_Cin(1);
			ELSIF (saida_deco(4)= '1') THEN
				S <= A_B_Cin(2) XOR A_B_Cin(1);
			ELSIF (saida_deco(5)= '1') THEN
				S <= A_B_Cin(2) XNOR A_B_Cin(1);
			ELSIF (saida_deco(6)= '1') THEN
				S <= S_Cout(1);
				Cout <= S_Cout(0);
			ELSIF (saida_deco(7)= '1') THEN
				S <= S_Cout2(1);
				Cout <= S_Cout2(0);
			END IF;		
		END PROCESS;
END COMPORTAMENTAL;