LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
		
COMPONENT NOT_1 IS
	PORT(A: IN BIT;
		 S: OUT BIT);
END COMPONENT;

COMPONENT AND_2 IS
	PORT(A,B: IN BIT;
		 S: OUT BIT);
END COMPONENT;

  
ENTITY DECODIFICADOR IS
	PORT(D0: IN BIT_VECTOR (1 DOWNTO 0);
		 SD0, SD1, SD2, SD3: OUT BIT_VECTOR (0 DOWNTO 0));
END DECODIFICADOR;

ARCHITECTURE TEST_DC OF DECODIFICADOR IS 
	BEGIN
		PROCESS (D0)
		BEGIN	
			CASE D0 IS
				WHEN "00" => SD0 <= "1" ;
				WHEN "01" => SD1 <= "1";
				WHEN "10" => SD2 <= "1";
				WHEN "11" => SD3 <= "1";
			END CASE;
		END PROCESS;
	END TEST_DC;
END DECODIFICADOR_PACKAGE;