LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CONT_SEG IS
	PORT(CLK, RST: IN BIT;
	     RCO: OUT BIT;
	     UNID, DEZ: OUT INTEGER RANGE 0 TO 15);
END CONT_SEG;

ARCHITECTURE COMPORTAMENTAL OF CONT_SEG IS 
	SIGNAL I0: BIT;
BEGIN
	UNIDADE: PROCESS(CLK,RST)
		VARIABLE CONT: INTEGER RANGE 0 TO 15;
	BEGIN
		IF (RST='0') THEN
			CONT:=0; I0 <='0';
		ELSIF (FALLING_EDGE(CLK)) THEN
			IF (CONT <9) THEN
				CONT:= CONT+1;
				CASE CONT IS
					WHEN 9 => I0 <='1'; WHEN OTHERS => I0 <='0';
				END CASE;
			ELSE CONT:=0; I0<='0';
			END IF;
		END IF;
		UNID<= CONT; -- UNIDADE ATUALIZADA
	END PROCESS UNIDADE;
	DEZENA: PROCESS(I0,RST)
		VARIABLE CONT: INTEGER RANGE 0 TO 15;
	BEGIN
		IF (RST='0') THEN
			CONT:=0; RCO <='0';
		ELSIF (FALLING_EDGE(CLK)) THEN
			IF (CONT<5) THEN
			CONT:= CONT +1;
			CASE CONT IS
				WHEN 5 => RCO <= '1'; WHEN OTHERS => RCO <='0';
			END CASE;
		ELSE CONT:=0; RCO <= '0';
		END IF;
	END IF;
		DEZ <= CONT; --DEZENAS ATUALIZADAS
	END PROCESS DEZENA;
END COMPORTAMENTAL;	
	
	     