-- SOMADOR COMPLETO DE 1 BIT
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SOMADOR IS
	PORT(A_B_Cin: IN BIT_VECTOR (2 DOWNTO 0);
		 S, Cout: OUT BIT_VECTOR (2 DOWNTO 0)); -- DA UMA VERIFICADA AQUI MAS ACHO QUE � S� 1 BIT QUE SAI
END SOMADOR;

-- O SOMADOR DEVE SER FEITO USANDO WHITE SELECT WHEN

ARCHITECTURE TEST_SOMADOR OF SOMADOR IS
	BEGIN
		WITH A_B_Cin SELECT
			S <= "0" WHEN "000" | "101" | "110" | "111",
			S <= "1" WHEN "001" | "010" | "100",
			Cout <= "0" WHEN "000",
			CouT <= "1" WHEN "010" | "001" | "100" | "111";
END TEST_SOMADOR;