LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
	
	-- DECLARA��O DOS COMPONENTES QUE IR�O COMPOR O MUX 2X1
	
--	COMPONENT AND_2 IS
--		PORT(A,B: IN BIT;
--			 S: OUT BIT);
--	END COMPONENT;
	
--	COMPONENT NOT_1 IS
--		PORT(A: IN BIT;
--			 S: OUT BIT);
--	COMPONENT NOT_1;
	
--	COMPONENT OR_2 IS
--		PORT(A,B: IN BIT;
--			 S: OUT BIT);
--	END COMPONENT;
	
	-- FIM DOS COMPONENTES
	-- INICIO DA ENTIDADE PARA O MUX 2X1
	
ENTITY MUX_2X1 IS
	PORT(A,B: IN BIT;
	     SEL: IN BIT; -- SELETOR DO MUX
		 Y: OUT BIT);
END MUX_2X1;

ARCHITECTURE TEST_MUX OF MUX_2X1 IS
	BEGIN
		PROCESS(A,B)
			BEGIN
				IF SEL = '0' THEN
					Y <= A AND NOT SEL;
				ELSE
					Y <= B AND SEL;
				END IF;
		END PROCESS;
	END TEST_MUX;
	