LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECODIFICADOR_8x1 IS
	PORT(E0,E1,E2,E3,E4,E5,E6,E7: IN BIT;
		 SAIDA_ULA: OUT BIT;
		 SEL: BIT_VECTOR (2 DOWNTO 0));
END DECODIFICADOR_8x1;

ARCHITECTURE TEST_DECO OF DECODIFICADOR_8x1 IS
BEGIN
	PROCESS(SEL,E1,E2,E3,E4,E5,E6,E7,E0)
		BEGIN
			CASE SEL IS
				WHEN "000" => SAIDA_ULA <= E0;
				WHEN "001" => SAIDA_ULA <= E1;
				WHEN "010" => SAIDA_ULA <= E2;
				WHEN "011" => SAIDA_ULA <= E3;
				WHEN "100" => SAIDA_ULA <= E4;
				WHEN "101" => SAIDA_ULA <= E5;
				WHEN "110" => SAIDA_ULA <= E6;
				WHEN "111" => SAIDA_ULA <= E7;
		END CASE;
	END PROCESS;
END TEST_DECO;

