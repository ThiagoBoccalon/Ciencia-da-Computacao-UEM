LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

	PACKAGE PORTAS_LOGICAS_PACKAGE IS
	
		COMPONENT NOT_1 IS
			PORT(A: IN BIT;
				 S: OUT BIT);
		END COMPONENT;
		
		COMPONENT AND_2 IS
			PORT(A,B: IN BIT;
				 S: OUT BIT);
		END COMPONENT;
		
		COMPONENT XOR_2 IS
			PORT(A,B: IN BIT;
				 S: OUT BIT);
		END COMPONENT;
		
	END PORTAS_LOGICAS_PACKAGE;
	
ENTITY PORTAS_LOGICAS IS
	PORT(E1, E2: IN BIT;
		 S1,S2: OUT BIT; -- S1 E S2 S�O SA�DAS PARA A UNIDADE L�GICA DA ULA.
		 S3,S4,S5,S6: OUT BIT);
END PORTAS_LOGICAS;

ARCHITECTURE TESTE_PORTA_LOGICAS OF PORTAS_LOGICAS IS
BEGIN
	PROCESS (E1, E2)
	BEGIN
		IF E1=E2 THEN
			S1 <= '1'; -- XNOR
			S2 <= '0'; -- XOR
		ELSE
			S1 <= '0'; -- XNOR
			S2 <= '1'; -- XOR
		END IF;
		
		IF E1='1' OR E2='1' THEN 
			S3 <= '0'; -- NOR
			S4 <= '1'; -- OR
		ELSE
			S3 <= '1'; -- NOR
			S4 <= '0'; -- OR
		END IF;
		
		IF E1='1' AND E2='1' THEN 
			S5 <= '0'; -- NAND
			S6 <= '1';  -- AND
		ELSE
			S5 <= '1'; -- NAND
			S6 <= '0';  -- AND
		END IF;
	END PROCESS;
END TESTE_PORTA_LOGICAS;
	