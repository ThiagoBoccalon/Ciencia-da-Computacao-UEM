library ieee;
use ieee.std_logic_1164.all;
entity Somador_1 is 
port (
generic ()
		);

architecture 