LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CONT_SINC_MOD4_C IS
	PORT(CLR,CLK: IN STD_LOGIC;
		 Q, QBAR: OUT )