LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY EXERCICIO_1_SELECT_WHEN IS
	PORT(CH: IN BIT_VECTOR(3 DOWNTO 0);
	     S: OUT BIT_VECTOR (3 DOWNTO 0));
END EXERCICIO_1_SELECT_WHEN;

ARCHITECTURE TEST_BETA OF EXERCICIO_1_SELECT_WHEN IS
BEGIN
		WITH CH SELECT
			S <= "0000" WHEN "0000",
			     "0001" WHEN "0001", -- DETALHE A VIRGULA
			     "0010" WHEN "0010" | "0011",
			     "0100" WHEN "0100" | "0101" | "0110" | "0111",
			     "1000" WHEN "1000" | "1001" | "1010" | "1011" | "1100" | "1101" | "1110" | "1111";
			     
END TEST_BETA;
			  
		