LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECODIFICADOR_3x8 IS 
	PORT(SEL: BIT_VECTOR (2 DOWNTO 0);
	--	 S : OUT BIT_VECTOR(7 DOWNTO 0));
		 S0,S1,S2,S3,S4,S5,S6,S7: OUT BIT_VECTOR (0 DOWNTO 0));
END DECODIFICADOR_3x8;

ARCHITECTURE TEST_DECO_3x8 OF DECODIFICADOR_3x8 IS
	BEGIN
		PROCESS(SEL)
			BEGIN
				CASE SEL IS
					WHEN "000" => S0 <= "1"; 
					WHEN "001" => S1 <= "1";
					WHEN "010" => S2 <= "1";
					WHEN "011" => S3 <= "1";
					WHEN "100" => S4 <= "1";
					WHEN "101" => S5 <= "1";
					WHEN "110" => S6 <= "1"; 
					WHEN "111" => S7 <= "1"; 
				END CASE;
			END PROCESS;
	END TEST_DECO_3x8;
		