LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY LATCH_D_CLK IS
	PORT(D, CLK: IN BIT; 
		 Q, QBAR: BUFFER BIT);
END LATCH_D_CLK;

ARCHITECTURE TEST_D_CLK OF LATCH_D_CLK IS
	BEGIN
		PROCESS(D,CLK)
			BEGIN
				IF (CLK = '1') THEN Q <= D; QBAR <= NOT D;
				ELSE Q <= Q; QBAR <= QBAR;
				END IF;
			END PROCESS;
		END TEST_D_CLK;
	