LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CONT_ASSIC_MOD4 IS
	PORT(CLR, CLK, ES: IN STD_LOGIC;
		Q_OUT, QB_OUT: BUFFER STD_LOGIC_VECTOR (1 DOWNTO 0));
END CONT_ASSIC_MOD4;

ARCHITECTURE ESTRUTURAL OF CONT_ASSIC_MOD4 IS

	COMPONENT FFT_C IS
		PORT(CLR, CLK, T: STD_LOGIC;
			 Q, QBAR: BUFFER STD_LOGIC);
	END COMPONENT;
	
BEGIN
	FFT_C1: FFT_C PORT MAP (CLR, CLK, ES, Q_OUT(1), QB_OUT(1));
	FFT_C2: FFT_C PORT MAP (CLR, Q_OUT(1), ES, Q_OUT(0), QB_OUT(0));
END ESTRUTURAL;