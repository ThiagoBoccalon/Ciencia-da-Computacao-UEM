LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FFT_C IS
	PORT(CLR, CLK, T: STD_LOGIC;
		 Q, QBAR: BUFFER STD_LOGIC);
END FFT_C;

ARCHITECTURE TESTE OF FFT_C IS
BEGIN
	PROCESS (CLR, CLK, T)
		VARIABLE QV, QBARV: STD_LOGIC;
	BEGIN
		IF (CLR = '0') THEN
			QV:= '0';
			QBARV:= NOT QV;
		ELSIF (FALLING_EDGE (CLK)) THEN
			IF (T ='1') THEN
				QV:=  NOT QV;
				QBARV:= NOT QV;
			ELSE
				QV:= QV;
				QBARV:= QBARV;
			END IF;
		END IF;
	Q<= QV; QBAR<= QBARV;
	END PROCESS;
END TESTE;