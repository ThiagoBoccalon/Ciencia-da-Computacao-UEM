LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY CONT_MOD4_EX1 IS
	PORT(CLR, CLK: IN BIT;
			Q: OUT INTEGER RANGE 0 TO 3);
END CONT_MOD4_EX1;

ARCHITECTURE COMPORTAMENTAL OF CONT_MOD4_EX1 IS
BEGIN
	PROCESS(CLR,CLK)
	VARIABLE CONT: INTEGER RANGE 0 TO 3;
		BEGIN
			IF (CLR='0') THEN
				CONT:=0;
			ELSIF(CLK'EVENT AND CLK='0') THEN
				IF (CONT < 3) THEN
					CONT:= CONT + 1;
					ELSE
						CONT:= 0;
				END IF;
			END IF;
			Q<= CONT;
	END PROCESS;
END COMPORTAMENTAL;