LIBRARY WORKTRABALHO;
USE WORKTRABALHO.blocos_package.all;
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY ULA IS
	PORT(A_B_Cin, SEL_ULA : IN BIT_VECTOR (2 DOWNTO 0);
		 --SAIDA_DECO: out BIT_VECTOR (7 DOWNTO 0);
		 --S_Cout,S_Cout2: out BIT_VECTOR(1 DOWNTO 0);
		 S, Cout : OUT BIT);
END ULA;
ARCHITECTURE TEST_ULA OF ULA IS
Signal t0,t1 : bit_vector(1 downto 0);
signal t3 : bit_vector (7 downto 0);
BEGIN
	P1: SOMADOR PORT MAP (A_B_Cin,t0);
	P2: SUBTRATOR PORT MAP (A_B_Cin,t1);
	P3: DECODIFICADOR_3X8 PORT MAP (SEL_ULA, t3);
	P4: PORTAS_LOGICAS PORT MAP(A_B_Cin,t3,t0,t1,S,Cout);
END TEST_ULA;
	