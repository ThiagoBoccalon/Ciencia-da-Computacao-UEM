LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REG_DESL IS
	PORT(CLR, CLK, SHIFTIN: IN STD_LOGIC;
	      SHIFTOUT: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END REG_DESL; -- SHIFTIN CORRESPONDE A ES SHIFTOUT CORRESPONDE A Qi

ARCHITECTURE COMPORTAMENTAL OF REG_DESL IS
SIGNAL SHIFT_BIT : STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN
	PROCESS(CLR,CLK,SHIFTIN)	
	BEGIN
		IF (CLR ='0') THEN
			SHIFT_BIT <= "0000";
		
		ELSIF (RISING_EDGE(CLK)) THEN
		--	IF (SHIFTIN='0') THEN
				SHIFT_BIT(3)<= SHIFTIN;
				SHIFT_BIT(2)<= SHIFT_BIT(3);
				SHIFT_BIT(1)<= SHIFT_BIT(2);
				SHIFT_BIT(0)<= SHIFT_BIT(1);
			END IF;
	--	END IF;
		END PROCESS;
		
		SHIFTOUT(3)<= SHIFT_BIT(3);
		SHIFTOUT(2)<= SHIFT_BIT(2);
		SHIFTOUT(1)<= SHIFT_BIT(1);
		SHIFTOUT(0)<= SHIFT_BIT(0);
END COMPORTAMENTAL;				