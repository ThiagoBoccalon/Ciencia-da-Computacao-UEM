LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE MUX_2X1_PACKAGE IS

COMPONENT NOT_1 IS
	PORT ( A: IN BIT;
           
			);
