LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY OR_3 IS  
	PORT(A,B,C: IN BIT;
		 S: OUT BIT);
END OR_3;

ARCHITECTURE TEST_4 OF OR_3 IS
BEGIN
	S <= A OR B OR C;
END TEST_4;