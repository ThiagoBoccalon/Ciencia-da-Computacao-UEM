LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY EXERCICIO_9_DEMUX_1X4 IS 
	PORT(A,B, E0: IN BIT;
		 S1,S2,S3,S4: OUT BIT);
END EXERCICIO_9_DEMUX_1X4;

ARCHITECTURE FLUXO_DE_DADOS OF EXERCICIO_9_DEMUX_1X4 IS
BEGIN	
	PROCESS (A,B,E0)
	BEGIN
		IF A='0' AND B='0' AND E0 ='1' THEN
					S1<= E0;
		ELSE
			IF A='1' AND B='0' THEN
					S2 <= E0;
			ELSE
				IF A='0' AND B='1' THEN
					S3 <= E0;
			     ELSE
					S4 <= E0;
				END IF;
			END IF;
		END IF;
	END	PROCESS;
END FLUXO_DE_DADOS;
		   	