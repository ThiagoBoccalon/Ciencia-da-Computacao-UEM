LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

	COMPONENT DECODIFICADOR_3x8 IS
		PORT (SEL: BIT_VECTOR (2 DOWNTO 0);
			  SAIDA_ULA: OUT BIT);
	END COMPONENT;
	
	COMPONENT DECODIFICADOR_8x1 IS
		PORT (SEL: BIT_VECTOR (2 DOWNTO 0);
			  E_SOM, E_SUB, E3, E4, E5, E6, E7, E8: IN BIT;	
			  SAIDA_ULA: OUT BIT);
	END COMPONENT;
	
	COMPONENT PORTAS_LOGICAS IS 
		PORT (A,B: IN BIT; -- AS PORTAs TER� 8 ENTRADAS AO TODO
			  ENT_PL: BIT_VECTOR (5 DOWNTO 0);
			  SAIDAS: BIT_VECTOR (5 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT SOMADOR IS
		PORT (A_B_Cin: IN BIT_VECTOR (2 DOWNTO 0);
			  S, Cout: OUT BIT_VECTOR (2 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT SUBTRATOR IS 
		PORT (EN_SUB: IN BIT_VECTOR (2 DOWNTO 0);
			  S_Cout: OUT BIT_VECTOR (1 DOWNTO 0));
	END COMPONENT;
	
	ENTITY ULA_1BIT IS
		PORT(
			 );
	
	ARCHITECTURE TEST_ULA OF ULA_1BIT IS
			SIGNAL 
		BEGIN
			
		
	