LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FLIPFLOPJK IS
	PORT(CLK, J,K: IN STD_LOGIC;
		 Q, QBAR: BUFFER STD_LOGIC);
END FLIPFLOPJK;

ARCHITECTURE TEST_JK OF FLIPFLOPJK IS
	BEGIN
		PROCESS(CLK,J,K)
			VARIABLE QV, QBARV: STD_LOGIC; -- BIT
			BEGIN
				IF (FALLING_EDGE(CLK)) THEN
					IF (J = '1' AND K = '0') THEN QV := '1'; QBARV := NOT QV;	
					ELSIF (J ='0' AND K='1') THEN QV:= '0'; QBARV := NOT QV;
					ELSIF (J = '1' AND K='1') THEN QV:= NOT QV; QBARV := NOT QV;
					ELSE QV:= QV; QBARV:= NOT QV;   -- ESSA VARIAVEL N�O PRECISA SER INICIALIZADA????
					END IF;
				END IF;
			Q<= QV; QBAR <= QBARV;
		END PROCESS;
	END TEST_JK;