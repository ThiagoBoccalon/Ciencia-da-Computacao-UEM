LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY AND_2 IS
	PORT(A,B: IN BIT;
		 S: OUT BIT);
END AND_2;

ARCHITECTURE TEST_1 OF AND_2 IS
BEGIN
	S <= A AND B;
END TEST_1;
