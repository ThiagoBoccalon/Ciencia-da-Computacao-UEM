LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY REG_DEL_EST IS
	PORT(CLR, CLK, ES: IN STD_LOGIC;
		 Q_OUT, QB_OUT: BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0));
END REG_DEL_EST;

ARCHITECTURE ESTRUTURAL OF REG_DEL_EST IS

COMPONENT FFD_C IS
	PORT(CLR, CLK, D: IN STD_LOGIC;
		 Q, QBAR: BUFFER STD_LOGIC);
END COMPONENT;

BEGIN
		FFD_C1: FFD_C PORT MAP (CLR,CLK,ES,Q_OUT(1),QB_OUT(1));
		FFD_C0: FFD_C PORT MAP (CLR,CLK,Q_OUT(1),Q_OUT(0),QB_OUT(0));
END ESTRUTURAL;		