LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY FLIPFLOPJK_CLRPST IS
	PORT(PST, CLR, CLK, J, K: IN STD_LOGIC;
		 Q, QBAR: BUFFER STD_LOGIC);
END FLIPFLOPJK_CLRPST;

ARCHITECTURE COMPORTAMENTAL OF FLIPFLOPJK_CLRPST IS
BEGIN
	PROCESS(PST, CLR)