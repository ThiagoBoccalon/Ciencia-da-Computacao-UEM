Library ieee;
Use ieee.std_logic_1164.all;
Package blocos_package is
COMPONENT PORTAS_LOGICAS IS
	PORT(A_B_Cin : IN BIT_VECTOR (2 DOWNTO 0);
		Saida_deco : IN BIT_VECTOR (7 DOWNTO 0);
		S_Cout, S_Cout2 : IN BIT_VECTOR (1 DOWNTO 0);
		S, Cout: OUT BIT);
END COMPONENT;
COMPONENT SOMADOR IS
	PORT (A_B_Cin: IN BIT_VECTOR (2 DOWNTO 0);    
		  S_Cout: OUT BIT_vector (1 DOWNTO 0));
END COMPONENT;

COMPONENT SUBTRATOR IS
	PORT(EN_SUB: IN BIT_VECTOR (2 DOWNTO 0);
		 S_Cout: OUT BIT_VECTOR (1 DOWNTO 0));
END COMPONENT;

COMPONENT DECODIFICADOR_3X8 IS
	PORT(SEL: BIT_VECTOR (2 DOWNTO 0);
		 S : OUT BIT_VECTOR(7 DOWNTO 0));
END COMPONENT;
end blocos_package;